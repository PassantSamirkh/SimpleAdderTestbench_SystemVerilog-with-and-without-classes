package adder_package;
	`include "driver.sv"
	`include "monitor_output.sv"
	`include "monitor_input.sv"
	`include "adder_checker.sv"
endpackage
	